// userInput module take in two button signals and 
module Input (clk, reset, KEYS, D);
	input logic clk, reset, KEYS;
	output logic D;
	Press up (.clk, .reset, .inputButton(KEYS) , .out(D));
	
	
endmodule

module Input_testbench();
	logic clk, reset, KEYS;
	logic D;
		
	// Set up the clock
	parameter CLOCK_PERIOD=100;
	initial begin
		clk <= 0;
		forever #(CLOCK_PERIOD/2) clk <= ~clk;
	end
	 
	Input dut (clk, reset, KEYS, D); 


	
	initial begin	
			reset <= 1;	 KEYS <= 0;			@(posedge clk);
													@(posedge clk); 
			reset <= 0; 					 @(posedge clk);
												 @(posedge clk);
												 @(posedge clk);
			KEYS <= 1;						 @(posedge clk);
													@(posedge clk);
										     	 @(posedge clk);
												@(posedge clk);
			reset <= 1;  KEYS<= 0; 	 	 @(posedge clk);
												 @(posedge clk);
												@(posedge clk);
												@(posedge clk);
			KEYS <= 1; 				 		@(posedge clk);
											@(posedge clk);
			reset<=1; 					@(posedge clk);
											@(posedge clk);
			
								
	$stop;
	end

endmodule